module ascii_convert
(
	input 
);






endmodule
